module ALU(
	input wire [1:0] ALU_Op;
	input wire [7:0] inA;
	input wire [7:0] inB;
	output reg isZero;
	output reg [7:0] out;
);

endmodule;
