module controller_tb;
reg clk;


endmodule
